package core_pkg;

  PTR_WIDTH = 32;
  
  INST_MEM_ADDR_WIDTH = 12;
  DATA_MEM_ADDR_WIDTH = 12;

endpackage
