package core_pkg;

  localparam DATA_WIDTH = 32;

  localparam INST_MEM_ADDR_WIDTH = 12;
  localparam DATA_MEM_ADDR_WIDTH = 12;

endpackage
